module combLogic(
  input w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008,
  output OscFlag // 输出震荡检测信号
);

  wire w_000_001, w_000_002, w_000_003, w_000_004, w_000_005;
  wire w_001_006, w_001_007, w_001_008, w_001_009, w_001_010;
  wire w_002_012, w_002_013, w_002_014, w_002_015;
  wire w_002_012_prev;  // 用于检测震荡的反馈信号

  // 原始逻辑电路（加入检测信号）
  not1    I001_001(w_000_001, w_000_002);
  and2    I001_002(w_000_002, w_003_001, w_000_003);
  and2    I001_003(w_000_004, w_003_002, w_000_005);
  and2    I001_004(w_001_006, w_000_005, w_003_003);
  and2    I001_005(w_001_007, w_003_004, w_000_003);
  and2    I001_006(w_001_008, w_000_001, w_000_004);
  nand2   I001_007(w_000_005, w_001_009, w_001_010);
  and2    I001_008(w_002_012, w_001_006, w_001_007);
  nand2   I001_009(w_000_003, w_002_013, w_002_014);
  nand2   I001_010(w_001_009, w_003_005, w_001_008);
  and2    I002_012(w_001_010, w_002_012_prev, w_003_006);
  and2    I002_013(w_002_013, w_003_007, w_002_012_prev);
  not1    I002_014(w_002_014, w_002_015);
  and2    I002_015(w_002_015, w_001_008, w_003_008);

  // 震荡检测逻辑
  // 定义一个简单的计数器计数 w_002_012 的变化次数
  wire change_detected = w_002_012 ^ w_002_012_prev;  // 检测w_002_012的状态变化
  wire [1:0] change_count;  // 用于记录变化次数

  // 组合逻辑版本的变化计数
  assign change_count = {w_002_012_prev, w_002_012} == 2'b01 ? 2 : 
                        {w_002_012_prev, w_002_012} == 2'b10 ? 2 : 1;

  // 当变化次数达到2次以上认为发生震荡
  assign OscFlag = (change_count >= 2) ? 1'b1 : 1'b0;

  // 反馈信号，用于保持电路在稳定态
  assign w_002_012_prev = w_002_012;

initial begin
    $monitor("Time=%t, OscFlag=%b", $time, OscFlag);
end

endmodule
