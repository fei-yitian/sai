module combLogic(w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, OscFlag);

  input w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008;
  output OscFlag;
  wire OscFlag;

  wire w_000_001, w_000_002, w_000_003, w_000_004, w_000_005;
  wire w_001_006, w_001_007, w_001_008, w_001_009, w_001_010;
  wire w_002_012, w_002_013, w_002_014, w_002_015;
  wire w_002_012_prev;  // 引入用于反馈控制的信号

  // 使用组合逻辑将 w_002_012 的上一状态反馈
  assign w_002_012_prev = w_002_012;

  not1    I001_001(w_000_001, w_000_002);
  and2    I001_002(w_000_002, w_003_001, w_000_003);
  and2    I001_003(w_000_004, w_003_002, w_000_005);
  and2    I001_004(w_001_006, w_000_005, w_003_003);
  and2    I001_005(w_001_007, w_003_004, w_000_003);
  and2    I001_006(w_001_008, w_000_001, w_000_004);
  nand2   I001_007(w_000_005, w_001_009, w_001_010);
  and2    I001_008(w_002_012, w_001_006, w_001_007);  
  nand2   I001_009(w_000_003, w_002_013, w_002_014);
  nand2   I001_010(w_001_009, w_003_005, w_001_008);
  and2    I002_012(w_001_010, w_002_012_prev, w_003_006);  // 使用 w_002_012_prev 控制反馈
  and2    I002_013(w_002_013, w_003_007, w_002_012_prev);
  not1    I002_014(w_002_014, w_002_015);
  and2    I002_015(w_002_015, w_001_008, w_003_008);

  // 检测震荡：如果 w_002_012 和 w_002_012_prev 的值频繁不同，则 OscFlag 为 1
  assign OscFlag = (w_002_012 != w_002_012_prev);

  initial begin
    $monitor("Time=%t, OscFlag=%b", $time, OscFlag);
  end
endmodule
